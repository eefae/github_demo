module test(){
};

endmodule
